`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.12.2023 18:17:11
// Design Name: 
// Module Name: tb_nexystop
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module tb_uartrx();
    reg CLK;
    reg RST;
    reg RX;
    
    uart_rx DUT(
        .clk_i(CLK),
        .rst_i(RST),
        .rx_i(RX)
    );
    initial CLK <= 0;
    always #50 CLK <= ~CLK;
    initial begin
        RST = 1;
        RX = 1;
        #100
        RST = 0;
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 1;
        
        #95680
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 0;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
        #8700
        RX = 1;
    end
    initial #3ms $finish();
    
endmodule
